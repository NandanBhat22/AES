module sTable(
  input [7:0] inByte,
  output reg [7:0] outByte
);


	always @(inByte) begin
		case (inByte)
			8'h00: outByte=8'h63;
			8'h01: outByte=8'h7c;
			8'h02: outByte=8'h77;
			8'h03: outByte=8'h7b;
			8'h04: outByte=8'hf2;
			8'h05: outByte=8'h6b;
			8'h06: outByte=8'h6f;
			8'h07: outByte=8'hc5;
			8'h08: outByte=8'h30;
			8'h09: outByte=8'h01;
			8'h0a: outByte=8'h67;
			8'h0b: outByte=8'h2b;
			8'h0c: outByte=8'hfe;
			8'h0d: outByte=8'hd7;
			8'h0e: outByte=8'hab;
			8'h0f: outByte=8'h76;
			8'h10: outByte=8'hca;
			8'h11: outByte=8'h82;
			8'h12: outByte=8'hc9;
			8'h13: outByte=8'h7d;
			8'h14: outByte=8'hfa;
			8'h15: outByte=8'h59;
			8'h16: outByte=8'h47;
			8'h17: outByte=8'hf0;
			8'h18: outByte=8'had;
			8'h19: outByte=8'hd4;
			8'h1a: outByte=8'ha2;
			8'h1b: outByte=8'haf;
			8'h1c: outByte=8'h9c;
			8'h1d: outByte=8'ha4;
			8'h1e: outByte=8'h72;
			8'h1f: outByte=8'hc0;
			8'h20: outByte=8'hb7;
			8'h21: outByte=8'hfd;
			8'h22: outByte=8'h93;
			8'h23: outByte=8'h26;
			8'h24: outByte=8'h36;
			8'h25: outByte=8'h3f;
			8'h26: outByte=8'hf7;
			8'h27: outByte=8'hcc;
			8'h28: outByte=8'h34;
			8'h29: outByte=8'ha5;
			8'h2a: outByte=8'he5;
			8'h2b: outByte=8'hf1;
			8'h2c: outByte=8'h71;
			8'h2d: outByte=8'hd8;
			8'h2e: outByte=8'h31;
			8'h2f: outByte=8'h15;
			8'h30: outByte=8'h04;
			8'h31: outByte=8'hc7;
			8'h32: outByte=8'h23;
			8'h33: outByte=8'hc3;
			8'h34: outByte=8'h18;
			8'h35: outByte=8'h96;
			8'h36: outByte=8'h05;
			8'h37: outByte=8'h9a;
			8'h38: outByte=8'h07;
			8'h39: outByte=8'h12;
			8'h3a: outByte=8'h80;
			8'h3b: outByte=8'he2;
			8'h3c: outByte=8'heb;
			8'h3d: outByte=8'h27;
			8'h3e: outByte=8'hb2;
			8'h3f: outByte=8'h75;
			8'h40: outByte=8'h09;
			8'h41: outByte=8'h83;
			8'h42: outByte=8'h2c;
			8'h43: outByte=8'h1a;
			8'h44: outByte=8'h1b;
			8'h45: outByte=8'h6e;
			8'h46: outByte=8'h5a;
			8'h47: outByte=8'ha0;
			8'h48: outByte=8'h52;
			8'h49: outByte=8'h3b;
			8'h4a: outByte=8'hd6;
			8'h4b: outByte=8'hb3;
			8'h4c: outByte=8'h29;
			8'h4d: outByte=8'he3;
			8'h4e: outByte=8'h2f;
			8'h4f: outByte=8'h84;
			8'h50: outByte=8'h53;
			8'h51: outByte=8'hd1;
			8'h52: outByte=8'h00;
			8'h53: outByte=8'hed;
			8'h54: outByte=8'h20;
			8'h55: outByte=8'hfc;
			8'h56: outByte=8'hb1;
			8'h57: outByte=8'h5b;
			8'h58: outByte=8'h6a;
			8'h59: outByte=8'hcb;
			8'h5a: outByte=8'hbe;
			8'h5b: outByte=8'h39;
			8'h5c: outByte=8'h4a;
			8'h5d: outByte=8'h4c;
			8'h5e: outByte=8'h58;
			8'h5f: outByte=8'hcf;
			8'h60: outByte=8'hd0;
			8'h61: outByte=8'hef;
			8'h62: outByte=8'haa;
			8'h63: outByte=8'hfb;
			8'h64: outByte=8'h43;
			8'h65: outByte=8'h4d;
			8'h66: outByte=8'h33;
			8'h67: outByte=8'h85;
			8'h68: outByte=8'h45;
			8'h69: outByte=8'hf9;
			8'h6a: outByte=8'h02;
			8'h6b: outByte=8'h7f;
			8'h6c: outByte=8'h50;
			8'h6d: outByte=8'h3c;
			8'h6e: outByte=8'h9f;
			8'h6f: outByte=8'ha8;
			8'h70: outByte=8'h51;
			8'h71: outByte=8'ha3;
			8'h72: outByte=8'h40;
			8'h73: outByte=8'h8f;
			8'h74: outByte=8'h92;
			8'h75: outByte=8'h9d;
			8'h76: outByte=8'h38;
			8'h77: outByte=8'hf5;
			8'h78: outByte=8'hbc;
			8'h79: outByte=8'hb6;
			8'h7a: outByte=8'hda;
			8'h7b: outByte=8'h21;
			8'h7c: outByte=8'h10;
			8'h7d: outByte=8'hff;
			8'h7e: outByte=8'hf3;
			8'h7f: outByte=8'hd2;
			8'h80: outByte=8'hcd;
			8'h81: outByte=8'h0c;
			8'h82: outByte=8'h13;
			8'h83: outByte=8'hec;
			8'h84: outByte=8'h5f;
			8'h85: outByte=8'h97;
			8'h86: outByte=8'h44;
			8'h87: outByte=8'h17;
			8'h88: outByte=8'hc4;
			8'h89: outByte=8'ha7;
			8'h8a: outByte=8'h7e;
			8'h8b: outByte=8'h3d;
			8'h8c: outByte=8'h64;
			8'h8d: outByte=8'h5d;
			8'h8e: outByte=8'h19;
			8'h8f: outByte=8'h73;
			8'h90: outByte=8'h60;
			8'h91: outByte=8'h81;
			8'h92: outByte=8'h4f;
			8'h93: outByte=8'hdc;
			8'h94: outByte=8'h22;
			8'h95: outByte=8'h2a;
			8'h96: outByte=8'h90;
			8'h97: outByte=8'h88;
			8'h98: outByte=8'h46;
			8'h99: outByte=8'hee;
			8'h9a: outByte=8'hb8;
			8'h9b: outByte=8'h14;
			8'h9c: outByte=8'hde;
			8'h9d: outByte=8'h5e;
			8'h9e: outByte=8'h0b;
			8'h9f: outByte=8'hdb;
			8'ha0: outByte=8'he0;
			8'ha1: outByte=8'h32;
			8'ha2: outByte=8'h3a;
			8'ha3: outByte=8'h0a;
			8'ha4: outByte=8'h49;
			8'ha5: outByte=8'h06;
			8'ha6: outByte=8'h24;
			8'ha7: outByte=8'h5c;
			8'ha8: outByte=8'hc2;
			8'ha9: outByte=8'hd3;
			8'haa: outByte=8'hac;
			8'hab: outByte=8'h62;
			8'hac: outByte=8'h91;
			8'had: outByte=8'h95;
			8'hae: outByte=8'he4;
			8'haf: outByte=8'h79;
			8'hb0: outByte=8'he7;
			8'hb1: outByte=8'hc8;
			8'hb2: outByte=8'h37;
			8'hb3: outByte=8'h6d;
			8'hb4: outByte=8'h8d;
			8'hb5: outByte=8'hd5;
			8'hb6: outByte=8'h4e;
			8'hb7: outByte=8'ha9;
			8'hb8: outByte=8'h6c;
			8'hb9: outByte=8'h56;
			8'hba: outByte=8'hf4;
			8'hbb: outByte=8'hea;
			8'hbc: outByte=8'h65;
			8'hbd: outByte=8'h7a;
			8'hbe: outByte=8'hae;
			8'hbf: outByte=8'h08;
			8'hc0: outByte=8'hba;
			8'hc1: outByte=8'h78;
			8'hc2: outByte=8'h25;
			8'hc3: outByte=8'h2e;
			8'hc4: outByte=8'h1c;
			8'hc5: outByte=8'ha6;
			8'hc6: outByte=8'hb4;
			8'hc7: outByte=8'hc6;
			8'hc8: outByte=8'he8;
			8'hc9: outByte=8'hdd;
			8'hca: outByte=8'h74;
			8'hcb: outByte=8'h1f;
			8'hcc: outByte=8'h4b;
			8'hcd: outByte=8'hbd;
			8'hce: outByte=8'h8b;
			8'hcf: outByte=8'h8a;
			8'hd0: outByte=8'h70;
			8'hd1: outByte=8'h3e;
			8'hd2: outByte=8'hb5;
			8'hd3: outByte=8'h66;
			8'hd4: outByte=8'h48;
			8'hd5: outByte=8'h03;
			8'hd6: outByte=8'hf6;
			8'hd7: outByte=8'h0e;
			8'hd8: outByte=8'h61;
			8'hd9: outByte=8'h35;
			8'hda: outByte=8'h57;
			8'hdb: outByte=8'hb9;
			8'hdc: outByte=8'h86;
			8'hdd: outByte=8'hc1;
			8'hde: outByte=8'h1d;
			8'hdf: outByte=8'h9e;
			8'he0: outByte=8'he1;
			8'he1: outByte=8'hf8;
			8'he2: outByte=8'h98;
			8'he3: outByte=8'h11;
			8'he4: outByte=8'h69;
			8'he5: outByte=8'hd9;
			8'he6: outByte=8'h8e;
			8'he7: outByte=8'h94;
			8'he8: outByte=8'h9b;
			8'he9: outByte=8'h1e;
			8'hea: outByte=8'h87;
			8'heb: outByte=8'he9;
			8'hec: outByte=8'hce;
			8'hed: outByte=8'h55;
			8'hee: outByte=8'h28;
			8'hef: outByte=8'hdf;
			8'hf0: outByte=8'h8c;
			8'hf1: outByte=8'ha1;
			8'hf2: outByte=8'h89;
			8'hf3: outByte=8'h0d;
			8'hf4: outByte=8'hbf;
			8'hf5: outByte=8'he6;
			8'hf6: outByte=8'h42;
			8'hf7: outByte=8'h68;
			8'hf8: outByte=8'h41;
			8'hf9: outByte=8'h99;
			8'hfa: outByte=8'h2d;
			8'hfb: outByte=8'h0f;
			8'hfc: outByte=8'hb0;
			8'hfd: outByte=8'h54;
			8'hfe: outByte=8'hbb;
			8'hff: outByte=8'h16;
		endcase
	end
endmodule
